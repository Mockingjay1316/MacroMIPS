module thinkpad_sv();
Clock clk;

